library verilog;
use verilog.vl_types.all;
entity JKFLIPFLOPUSINGIFELSE_vlg_check_tst is
    port(
        q               : in     vl_logic;
        qb              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end JKFLIPFLOPUSINGIFELSE_vlg_check_tst;
