library verilog;
use verilog.vl_types.all;
entity JKFLIPFLOPUSINGIFELSE_vlg_vec_tst is
end JKFLIPFLOPUSINGIFELSE_vlg_vec_tst;
